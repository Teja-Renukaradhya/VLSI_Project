magic
tech scmos
timestamp 1460680199
<< nwell >>
rect -20 -2 -10 16
rect 7 -2 17 16
rect 46 11 66 21
rect 46 -34 69 -23
<< polysilicon >>
rect 55 36 96 38
rect -26 31 32 33
rect -26 8 -24 31
rect -26 6 -18 8
rect -12 6 -8 8
rect -3 6 9 8
rect 15 6 20 8
rect 30 7 32 31
rect 55 19 57 36
rect 55 8 57 13
rect -26 -26 -24 6
rect -3 -26 -1 6
rect 55 -6 57 -3
rect 26 -18 28 -12
rect 55 -18 57 -12
rect 26 -20 57 -18
rect 55 -26 57 -20
rect -26 -28 -18 -26
rect -12 -28 -8 -26
rect -3 -28 9 -26
rect 15 -28 20 -26
rect -3 -69 -1 -28
rect 55 -39 57 -31
rect 56 -58 58 -56
rect 56 -69 58 -64
rect 94 -69 96 36
rect -3 -71 96 -69
<< ndiffusion >>
rect -18 -24 -17 -20
rect -13 -24 -12 -20
rect -18 -26 -12 -24
rect 48 -10 49 -6
rect 53 -10 55 -6
rect 48 -12 55 -10
rect 57 -10 58 -6
rect 62 -10 63 -6
rect 57 -12 63 -10
rect 9 -23 10 -19
rect 14 -23 15 -19
rect 9 -26 15 -23
rect -18 -30 -12 -28
rect -18 -34 -17 -30
rect -13 -34 -12 -30
rect 9 -29 15 -28
rect 9 -33 10 -29
rect 14 -33 15 -29
rect 48 -62 50 -58
rect 54 -62 56 -58
rect 48 -64 56 -62
rect 58 -62 60 -58
rect 64 -62 66 -58
rect 58 -64 66 -62
<< pdiffusion >>
rect -18 10 -17 14
rect -13 10 -12 14
rect -18 8 -12 10
rect 9 10 10 14
rect 14 10 15 14
rect 9 8 15 10
rect 48 15 49 19
rect 53 15 55 19
rect 48 13 55 15
rect 57 15 58 19
rect 62 15 64 19
rect 57 13 64 15
rect -18 4 -12 6
rect -18 0 -17 4
rect -13 0 -12 4
rect 9 4 15 6
rect 9 0 10 4
rect 14 0 15 4
rect 48 -27 55 -26
rect 48 -31 50 -27
rect 54 -31 55 -27
rect 57 -27 67 -26
rect 57 -31 60 -27
rect 64 -31 67 -27
<< metal1 >>
rect -17 25 14 28
rect -17 14 -13 25
rect -9 21 3 25
rect 7 21 14 25
rect 10 14 14 21
rect 49 7 53 15
rect -17 -8 -13 0
rect -33 -12 -13 -8
rect -33 -76 -29 -12
rect -17 -20 -13 -12
rect 33 3 53 7
rect 10 -8 14 0
rect 49 -6 53 3
rect 10 -12 25 -8
rect 58 -6 62 15
rect 62 -10 85 -7
rect 10 -19 14 -12
rect 50 -27 54 -26
rect -17 -44 -13 -34
rect 10 -40 14 -33
rect -9 -44 3 -40
rect 7 -44 14 -40
rect 50 -58 54 -31
rect 60 -27 64 -26
rect 82 -27 85 -10
rect 64 -30 85 -27
rect 60 -58 64 -31
rect 50 -76 54 -62
rect -33 -80 54 -76
<< ntransistor >>
rect 55 -12 57 -6
rect -18 -28 -12 -26
rect 9 -28 15 -26
rect 56 -64 58 -58
<< ptransistor >>
rect -18 6 -12 8
rect 9 6 15 8
rect 55 13 57 19
rect 55 -31 57 -26
<< polycontact >>
rect 29 3 33 7
rect 25 -12 29 -8
<< ndcontact >>
rect -17 -24 -13 -20
rect 49 -10 53 -6
rect 58 -10 62 -6
rect 10 -23 14 -19
rect -17 -34 -13 -30
rect 10 -33 14 -29
rect 50 -62 54 -58
rect 60 -62 64 -58
<< pdcontact >>
rect -17 10 -13 14
rect 10 10 14 14
rect 49 15 53 19
rect 58 15 62 19
rect -17 0 -13 4
rect 10 0 14 4
rect 50 -31 54 -27
rect 60 -31 64 -27
<< psubstratepcontact >>
rect -13 -44 -9 -40
rect 3 -44 7 -40
<< nsubstratencontact >>
rect -13 21 -9 25
rect 3 21 7 25
<< labels >>
rlabel polysilicon -25 -4 -25 -4 1 A
rlabel polysilicon -2 -5 -2 -5 1 B
rlabel metal1 84 -18 84 -18 1 Vo
rlabel metal1 -5 -42 -5 -42 1 gnd
rlabel metal1 -3 27 -3 27 1 VDD
<< end >>
