* SPICE3 file created from xor1.ext - technology: scmos

.model pfet pmos
.model nfet nmos

.tran 0.05n 40n


M1000 VDD A a_n18_n26# w_n20_n2# pfet w=6u l=2u
+ ad=72p pd=48u as=71p ps=48u
M1001 VDD B a_9_n26# w_7_n2# pfet w=6u l=2u
+ ad=0p pd=0u as=36p ps=24u
M1002 Vo B A w_46_11# pfet w=6u l=2u
+ ad=92p pd=56u as=42p ps=26u
M1003 Vo a_9_n26# A Gnd nfet w=6u l=2u
+ ad=84p pd=52u as=42p ps=26u
M1004 a_n18_n26# A gnd Gnd nfet w=6u l=2u
+ ad=84p pd=52u as=66p ps=46u
M1005 a_9_n26# B gnd Gnd nfet w=6u l=2u
+ ad=42p pd=26u as=0p ps=0u
M1006 Vo a_9_n26# a_n18_n26# w_46_n34# pfet w=5u l=2u
+ ad=0p pd=0u as=0p ps=0u
M1007 Vo B a_n18_n26# Gnd nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u


C0 gnd gnd! 6.4fF
C1 a_9_n26# gnd! 20.3fF
C2 a_n18_n26# gnd! 40.8fF
C3 Vo gnd! 15.5fF
C4 VDD gnd! 10.6fF
C5 A gnd! 45.8fF
C6 B gnd! 89.7fF

VDD VDD 0 5
vgnd gnd! 0 0
VA A 0 0 pulse 0 5 5n 2n 2n 10n 20n
VB B 0 0 pulse 0 6.0 2n 2n 2n 5n 20n
.probe V(A) V(B) V(Vo)
.End
