magic
tech scmos
timestamp 1460672980
<< nwell >>
rect -21 9 24 21
<< polysilicon >>
rect -8 18 -6 23
rect 9 18 11 23
rect -8 -2 -6 12
rect -17 -4 -6 -2
rect -8 -21 -6 -4
rect 9 6 11 12
rect 9 4 20 6
rect 9 -21 11 4
rect -8 -30 -6 -27
rect 9 -30 11 -27
<< ndiffusion >>
rect -18 -23 -8 -21
rect -18 -27 -14 -23
rect -10 -27 -8 -23
rect -6 -27 9 -21
rect 11 -23 21 -21
rect 11 -27 15 -23
rect 19 -27 21 -23
<< pdiffusion >>
rect -18 14 -16 18
rect -12 14 -8 18
rect -18 12 -8 14
rect -6 14 -3 18
rect 1 14 9 18
rect -6 12 9 14
rect 11 14 15 18
rect 19 14 21 18
rect 11 12 21 14
<< metal1 >>
rect -18 31 -16 35
rect -12 31 -2 35
rect 2 31 15 35
rect 19 31 21 35
rect -16 18 -12 31
rect 15 18 19 31
rect -16 12 -12 14
rect -3 2 1 14
rect 15 12 19 14
rect -3 -2 19 2
rect 15 -7 19 -2
rect 15 -11 27 -7
rect 15 -23 19 -11
rect -14 -37 -10 -27
rect -18 -41 -14 -37
rect -10 -41 15 -37
rect 19 -41 21 -37
<< ntransistor >>
rect -8 -27 -6 -21
rect 9 -27 11 -21
<< ptransistor >>
rect -8 12 -6 18
rect 9 12 11 18
<< ndcontact >>
rect -14 -27 -10 -23
rect 15 -27 19 -23
<< pdcontact >>
rect -16 14 -12 18
rect -3 14 1 18
rect 15 14 19 18
<< psubstratepcontact >>
rect -14 -41 -10 -37
rect 15 -41 19 -37
<< nsubstratencontact >>
rect -16 31 -12 35
rect -2 31 2 35
rect 15 31 19 35
<< labels >>
rlabel metal1 23 -9 23 -9 7 vout
rlabel polysilicon -16 -3 -16 -3 3 A
rlabel polysilicon 16 5 16 5 1 B
rlabel metal1 6 33 6 33 5 VDD
rlabel metal1 1 -39 1 -39 1 gnd
<< end >>
